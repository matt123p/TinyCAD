library ieee;
use ieee.std_logic_1164.all;

entity SINK is
	port(I0: in std_logic);
end SINK;

architecture structural of SINK is

begin
end structural;

